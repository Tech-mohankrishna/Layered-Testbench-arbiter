interface intf(input logic clk);
  logic reset;
  logic d;
  logic q;
  logic qb;
  
endinterface